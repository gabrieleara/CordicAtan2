library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity System_TB is
end System_TB;

architecture System_TB_Arch of System_TB is

	component CORDICAtan2 is
		port (
			clock			: in	std_ulogic;
			reset			: in	std_ulogic;
			inA				: in	std_ulogic_vector(12-1 downto 0);
			inB				: in	std_ulogic_vector(12-1 downto 0);
			valid			: out	std_ulogic;
			atan2Out		: out	std_ulogic_vector(12-1 downto 0)
		);
	end component;

	constant SIZE			: positive := 12;
	constant LUT_SIZE		: positive := 11;
	constant TEST_SIZE		: positive := 1000;

	type word_array			is array (natural range <>) of
        std_ulogic_vector(SIZE-1 downto 0);

	signal test_inA			: std_ulogic_vector(SIZE-1 downto 0);
	signal test_inB			: std_ulogic_vector(SIZE-1 downto 0);
	signal test_output		: std_ulogic_vector(SIZE-1 downto 0);
	signal test_valid		: std_ulogic;

	signal test_expected	: std_ulogic_vector(SIZE-1 downto 0);

	signal test_correct		: std_ulogic := '1';
	signal test_reset		: std_ulogic := '1';
	signal test_clock		: std_ulogic := '0';
	signal test_end			: std_ulogic := '0';

	-- TODO: fill these
	constant test_inputA		: word_array := ("110001100111","000101111001","011101100100","111010110111","101000110101","010100010010","010001000010","001000011100","001011100110","111001100111","010000001101","010110100110","100011110110","101101110110","110100001000","101110000000","101010110110","101111111010","001101001000","101000011000","000111111001","101000100000","001010010101","111100010111","101100110011","001010100001","111101010010","100001000000","111101111101","010110010111","000100001110","001011011010","101000110110","101001011100","001100011011","110001011101","000011111111","011000101001","000101011010","100011000110","100111011001","000011111010","011111001010","100000101001","111000101010","000000011110","010010001010","011000000110","100110110001","110011111011","010101010001","011100010111","011100000111","101101011100","010001011101","010111110100","000111111000","011110011000","101010010011","001001111010","011001000111","111011110110","010011011000","011000110100","100100010011","110101100111","001011111001","100011101110","001101111110","100000001000","101000101000","010010101101","111011011100","001010110000","011010101101","011101010111","101010000011","011110111111","011110010001","010100011000","110100100110","100110111101","100001000010","100000000110","101001111010","011100000000","111000010011","001101100111","111100111110","000011000110","011111111110","101100001111","111101100010","101000100011","100100100111","111000101100","011011101011","001010100101","010000110101","011001100000","011010011110","011011111000","110011010111","101000001101","000011111110","100000101100","100111000011","000001101100","011101011110","111010011000","011001001000","100000110001","110011010110","010100000011","010110010110","001001001001","100100010001","011001110110","111011111000","011101111110","101000101100","000001100111","110001101110","110110001101","101111010010","101000110100","000010101001","001010011010","000010110110","100001101001","100101011101","010110000100","101100000011","010010110110","011010110001","100001000011","000110011101","001111100100","100101011111","001101010110","101001010101","100001111111","110011111010","000001111110","000010010101","101001000001","111101110001","010110110101","111010100100","111000101000","110101010111","011011100011","011001110001","110110101000","110111000010","011100001001","101010010100","010011010000","100010010101","110110100001","010101100011","111010110001","000001111000","000011100101","001000100010","100110001001","011000110111","011010001111","110000101011","001111000101","101001100100","001010011000","111010011001","101101011000","001111111011","100101100110","101111001001","000010010011","110100011110","000111001011","000001110000","001010000101","111010001111","110001110001","011100100010","111110011101","010011010010","001110001010","001010001001","001101101010","011001010111","101110100100","111010001101","110100101001","111001010111","000011111000","010100011010","011010110000","011001010011","000110010101","001110110001","010111100011","111010100010","001001110101","101101100111","001001101111","110011111110","101111010011","100010000100","011011010111","111100011010","011001110100","001010001011","011010100111","111011110100","011111101100","110101100110","100001101010","100101101111","011110100110","000011001110","111000001000","111001010001","111001000100","110011101010","101111001110","000111100110","011001110101","110110111011","100001111110","111100101110","100010110000","011010000101","100110110100","010001001100","011110111000","010001010011","101101110100","100101011000","111100001011","010000110100","011000110010","100110101101","110110101111","001011101001","101100100001","010101100000","011101111100","010110110000","100011010001","100001001101","011101111101","000111101111","100010111010","001011111011","000101101111","001010111000","110010000101","110101111001","001010000001","011000101000","000110110001","010101001110","001011011011","101010101100","110101001010","100011100011","100111100101","000111011111","110101001011","100111010101","101101111111","011110101111","110111001100","001110000101","100011111111","011101010000","101001000111","111000111011","000011101000","100001001000","000100010111","100010000010","101111001100","110000110111","110101011011","100110000010","010111110000","100001111000","111110001011","101111001111","110101111011","101011010010","011110010110","001000101000","001100101111","100110110000","100011000001","010111010011","100001001100","011011100001","000111110101","011000110110","001010110001","010010100000","100011010111","100010000110","010111101100","100000110110","001110110100","111011010100","111101011010","111110101101","110101101011","001100000010","110001011010","101100100010","100110110111","101110011100","100101110011","101010000101","100101111111","000101110101","100111111010","011100101011","001111101000","111100101101","001101001110","100100001111","111001001011","111011111110","101010110111","110101110001","111011110101","101001000000","100010101111","000100001111","100011011100","000000100110","111111000111","011101000001","100000110101","010000010000","100000110100","001011001000","111111111000","111000000001","111110011100","100011011011","000000111000","001100000000","111000100111","100010110011","101100011100","110010011101","100011000000","010110000010","010000100001","110001100100","010011000011","000100111001","110100000010","110000010011","101001101111","001001111000","100001110010","010100011111","001100111011","100111100010","101111001000","110010110001","000110001001","011000011011","011001000000","000011011111","101110000111","011110110101","001001001100","100100101011","100101010011","110000100110","011100101001","110001000111","010011101110","111101011101","110100110011","100101110100","001100110011","010011100110","101001011110","101110110101","100110110010","101111000000","100110010011","000010011000","011010100001","111011101110","000001000011","101001010000","010110111010","011000010010","111110100111","100000011001","111110010010","101110001110","000000000000","011100011000","101010100100","001101101111","101111110000","001111000110","010111011011","010110001101","010111111010","110011111001","000101001100","101111101110","110010011011","011000100011","111101000101","001001101101","010001011010","011001001110","111101110110","110000111101","000000111011","111110101010","001101110010","111011011001","100100011100","101011000101","110111110011","111001011000","100010000101","000000011100","000000011001","001111110100","100100100001","010000111110","010000000111","001100001001","001111011111","001011001001","111101111000","111111001100","000101010001","000001010111","000011010111","011011001010","110001110000","111001001111","110001010001","001101100101","100110101100","100010111001","111101001000","010000110001","011010001101","100000010111","100110010110","110011011001","010101001001","100011110001","101110100010","100100101010","000000110110","010101000111","110111000001","101111011000","000100000101","111000111110","101011111111","101110010010","010111101010","111100000011","110000010110","100100011111","101110010100","111110000100","110000100111","010110111101","111001111001","001010010010","011001110011","001111011010","011100111101","010101001000","011111100111","010110101010","010100100100","101101001110","011001111111","100100101100","101000000011","001110011110","011111110001","000001111111","110000001100","110001000100","101100001000","110110111110","100001001010","110001111111","001110001111","001111111101","000000101011","001000001111","001110100011","111001001001","100100111000","010110101100","100100010101","110010000010","011000101111","110110100010","011000101100","101000110010","101011110011","100011000010","101000111111","011110101000","101100011000","100101101010","110101110111","101001111100","001100110001","110111010101","101110000100","110111100010","011001100110","101101001111","101000100001","000011000111","000101010111","001010101110","100110010010","000000110011","001110010101","111100010101","111111101101","100110111010","111010111000","010110100111","101000000000","011011000001","101100011011","001101111101","101111010101","100111010010","011101110110","100001010000","011100100101","001011000110","000110001000","101010001011","111001001010","111101011011","101100111110","110111000100","000011101110","101010100110","111001010101","000110110101","011110011111","100111111100","001011001010","100010010010","010111011100","100001011010","001010110111","010100101011","011111001111","101000000010","001111000000","010111110101","011101100011","001100100101","101110000101","011101000110","000011000101","011000110011","111000000110","010010010111","110100011100","100011001101","010000010100","010110001100","000110011001","010101111111","011011111100","010000100000","000001110101","001100011001","100000011000","101010110000","010011001000","101001100010","000010011001","100100001001","101110010110","010000011000","100111000000","101011110100","110101000111","010011110010","011111100011","111101000000","111101100000","000101100000","100111001111","010010011101","101000100100","110010010001","110010110101","110101111010","101011010001","110100001010","111100011011","011000110001","000010110100","010001010000","011110110010","111000001100","011010001011","110101101010","010110100101","100011010101","100101011100","100101111001","101001100101","001001100110","101101000000","001100101011","011100111011","100101111011","011000100100","110101001110","010100010110","101000111000","000111110011","011000111101","011010101110","000110110000","100010100011","000001111100","111101000010","101101110111","100110001010","110101100101","001001000000","011100100011","011000100111","111100010000","010010010000","000110101101","101001110101","111011100000","111110110101","101010001100","010001111100","010101111011","000000000011","101001001110","000001001011","110101101111","101100110000","110011001000","100001101111","000110000001","011110100100","100101010010","110000101111","100111101001","110111111110","110110101101","001111111110","011000101110","011011010001","000010001011","000001010001","101011011000","110101101110","001010010110","010100011100","110101110000","100110101110","101100101101","111001110100","000000101101","011010100100","001000011001","101001110110","111110100001","010111001111","110100010100","011100101100","010000000101","011101110011","110001000001","110110010000","010000101100","101000110111","010101010010","101001011111","100100101101","100001110110","000001100110","101001000010","001000101101","010101110100","111001101110","011101101011","101000001100","011111001011","000001001110","101100001100","010111100010","000101111010","010001100001","110011100110","000100101101","110010011001","011111001001","111010010011","010100010100","010001100000","010001001010","100010010011","010100111110","111110011000","110011110110","111010101010","000010111011","110000000010","010110100000","000011010110","110011101001","110111100100","011101111010","110101000000","101111100111","100100100110","000110111011","001001111001","111001100001","001010000010","010101111000","000001100011","010101100010","001101111100","110001000011","001101101100","111111111010","000110100110","110011111000","010001000110","111110101000","100101100100","010010010110","010101101100","110110011011","101010101101","001011110110","000000001001","101001100110","110101111100","111100100001","110000010000","110011001110","110000100000","111100011000","100010000000","010010000101","101011011100","100111101110","010010111010","000000011101","011010010101","101010110001","111010000111","101110000001","011000110101","011111010101","010010000111","110101100000","011010100011","011101001000","111000101110","001111011100","101001000110","011001011101","001000000111","100111100011","101111101101","111011000000","100000101010","110000110101","011001100111","101000101010","011101000010","101011110001","111011110111","101110001101","101001011101","001111101010","110011010001","001110000100","000001011000","001001100011","111110101110","000011010100","000111110010","010100010101","110101001001","010011011111","100011001110","110000111000","101110101110","110101101000","111010100111","100100111101","011011001110","111000101011","001110011001","101111111011","001011100011","101111110001","011110010111","011100111000","001010101011","100101110101","110010010010","001001110000","111010001110","100011100111","101011011001","000100000001","010001001101","011011000000","100111011010","011001100011","001010111101","011110001111","100011011110","111001011100","011010111001","111010010110","000111001000","001101101110","010101101110","010000001110","010110010001","001000001100","001111110001","011111001100","000110000000","101001001011","111011101111","011000100001","011100100001","110100001110","110100100010","111110010100","101100001110","011111010110","110000010001","111101110011","010011111000","010001000111","010111110110","101011100010","100011101111","011110001011","111011011110","011011010101","011111010100","000101100100","110010111110","111010101001","001001000001","000101001010","001110110101","010000111111","011110100000","110001001011","000001001101","101101001101","001001111110","110001000000","100101100001","010111110111","010010101110","111010111001","100100000111","111010101110","100011101101","101011100101","011010010110","101001110010","101000011101","001001000110","011101001111","011000000011","000011101111","100110001000","110110000110","100110101000","100111011100","111101110101","010100001010","011111101110","100011000100","111010100000","011010110100","011010011000","110101010100","100000100000","101110001011","011011101110","011111000110","100001100001","000111010011","101110110011","110100000001","000110110111","000111111101","011111011011","011100100110","111010001001","101011000111","111110111110","000010011011","001111001110","010101111110","100010010001","000011001000","001001011100","000010000011","101010111001","101110111011","111111000000","110011100100","011011000110","000001001001","010111100100","001011110111","110111110010","011110010010","111111100001","111101000111","111010110010","100000001110","101010101010","101100110100","110110000001","100001001001","011011101111","010111110011","000000011000","110111011000","000001100101","010100100000","101101111001","011100110100","011000000000","001100101110","010100000110","011011110111","101110010101","000000000000","010101101101","111000000010","111100011111","011001001001","101010110100","100011000101","100000010101","110110001011","100001100000","111110001101","110100011010","011010111010","101110100001","110000110100","001110101010","111101100100","101111010100","001001101000","001101110100","101101111110","010011000101","001001011111","110011000001","111110110010","001001010000","011000001000","001001011000","011001100010","010111110010","110000010100");
	constant test_inputB		: word_array := ("001011110100","000111000000","000110110100","100110010100","010011000100","010111001010","111111011100","110010101100","110011010001","101110001101","110011011011","000101001010","011100000010","110110101100","001101011011","101101001110","011001010010","100110100001","100010011100","000101011000","101001010100","101111001011","011100010010","000101010010","110111000010","001111101010","001011000100","110101101111","001100110101","111110110000","011100000111","011011110001","101010000110","010001110111","011001100100","000100000101","010111111100","001001110101","110111010101","000001101010","010001110001","110011110101","100010001000","101001100010","110001110000","101001001111","010100000101","001001101010","001111110001","000001001111","100001101010","010000110000","111101011001","011000111001","001111101011","010111001101","001111110100","101101110011","101101000001","001000011100","000101110100","001101101010","001110110011","001010011110","100010101000","101001000000","100100011110","100000011010","110110101010","010100000010","011101111001","111000110111","001001000011","011001100010","000101110110","101101011100","001000110001","011111100011","101001111100","000001111000","011000001010","101000000111","101101001100","101010010110","001001010011","100100010101","000110001100","011110010100","000101110011","001011001110","011011011000","010000110110","001100110000","110000001100","111100001000","011101011101","011001011010","101111110110","010110100010","010110000000","011111101101","100000101001","001110111110","011100100011","100010111001","000101000000","000001001100","100011101011","010100001000","011110000100","101011000111","010101110100","111111010010","101100010011","000110101000","001110001010","011100010100","101000110111","100101001100","101110101110","110011101101","110010101000","110111100111","001110110100","100001101110","001010100000","110001000111","110000110001","000011100001","100110101101","101110111101","110010001001","110101001110","110111010010","000101011001","110011110000","001011110001","001110001111","111110001001","111000011100","011110110010","111001011101","000100100110","110010011111","111000111010","100011000001","010001101000","100100011001","010101001110","001011101011","100011110101","111000101000","010100001110","111001110010","111110101000","110011001111","011101101110","101100000001","010101101101","101000111000","011011000101","111010001101","111011100011","100100100010","011011011001","001010010111","010110101011","001000011000","111110010101","100011001100","111100111001","111110101011","110011010100","001111001011","101011101001","001111000100","010011010000","001100111101","011100111110","011010001111","101100111011","110101001000","110010111011","011010000011","000001001001","010100101001","001011000101","011010111101","011001011111","100011100110","000011101001","010111100101","010101110101","101101001111","101000011001","111001001101","111100010010","001000011110","011100011010","111011111011","011100101011","111000000111","111011000111","001001010010","010010011100","010001011101","100011011111","110101000001","000000011100","011001000111","111101010111","101011011111","100001110101","111111111001","010001110100","110001100000","100011010110","010011111001","001111001001","111100011110","001111000010","010100010101","011010110111","000000111101","101010011100","001011011000","101010111100","111000010000","111011100001","000000010011","000111011011","100000001000","011101110100","010011001110","100110001100","011110011111","100101110000","101110010100","110101110000","000111100101","000001011101","110101101100","011010110000","110101000000","110100010110","111000010100","110111000110","110000001000","110001100110","111101001010","011100011000","100110110001","111000101100","000000011011","101110100000","010001111100","101011101101","011001111010","111111001110","110111101011","100001110100","011100101000","110100011000","001111111100","000010000001","101011100001","000100101110","001010010010","011111011110","111111001001","100001100111","110010011000","101001011100","000001000100","110010111111","111001100010","111001011000","100101100101","101100100010","101110110010","100011010000","000101001000","101100010010","000001101110","111111010111","000011110101","000011111111","100111001000","010110111100","001100000101","011111101111","000001000011","001010001110","000011101111","100110001111","101000111010","110011110111","010101000000","100001011001","101011001100","110110110110","110001110010","111011110000","010000011010","001010111011","001011110011","110000101010","101001000011","111000110001","000110100100","011110110100","111010000100","000011110111","110110010001","010100101111","101010001110","110010001110","000010000111","111100101011","111011111010","010110001011","010101001000","100100001100","110100110011","101010010010","110010011010","100000000010","011101010001","110011110011","001100111011","110101011100","100100000000","101010011010","011110111110","100101001000","111001100110","110110101111","000100111111","010101100100","001001011010","011010010100","010101100110","000101000101","110101010011","000100001100","010001000100","111011000010","110010100111","111010111000","100111100001","100100110010","111010011101","111111101100","000000110000","010010110000","111100010000","101011111000","110000111010","101101111010","100010001110","011111111001","100000100001","011010010111","110100111100","011101110000","110001010110","110111001101","010100000000","000010000110","111001000110","001100110111","100010100011","011111011000","111010111001","001101110101","010111000101","000010011110","010000101111","101101100110","111011010101","000101000111","011100001001","101111000100","000011010111","001110000100","001001110110","100010000011","010110110100","101100001101","011111011010","110010111001","011101100100","011101010110","101011100100","001001010100","011001110011","100101101011","001101101110","010110000011","010010101000","100110100010","011110000011","100011110100","111010101010","100000011011","001100111001","011000011101","000101010101","011111110001","110111011100","010100110000","100101011000","110001011000","110101100111","011001001110","000000011010","100000000100","011000010001","010011100010","000011110100","100100011011","111000010101","101000100100","101100010001","001111101100","110010101101","101010100111","101111011111","000111110001","111111100111","100110011000","100011100100","100001001111","000001110010","011001000110","111111011000","011011001011","111001011010","100011110011","011001101111","110010010111","101000001010","000111000001","011110011000","110000100011","001000111001","100001000100","111111111000","000000001001","010001110011","000111000111","111000000000","010000101110","001010001010","010010110100","100101110101","100111111011","100001001011","000101101100","001100110001","110000011100","011011010110","011011111110","100101010111","100000010011","110011000100","111101111111","000001011000","110100010010","100111100010","001001011110","010011111010","101000011100","000110111101","000110100101","101000001110","111010000001","101001100111","100000011000","010101100101","001001101111","010011010011","001001011111","101111010110","010000100010","110011110010","010010011111","111100011101","000110110010","001110001011","001100011001","001110100000","111110010111","010010110110","011101110110","011101011001","001110000011","011011011010","000100111001","110100100010","000100111011","010110110001","000000000001","000111111111","100010110010","000110110011","000001111111","011111101100","110000011000","001001001101","000010001100","011000001110","101001010010","111000100111","000010101001","111010001000","010010001111","101000101110","001111110010","000110110111","100111010011","111101000100","101101100010","011010001110","001110101110","110110010110","111111000001","100101010100","100001000111","010100011011","111011011100","000110100010","010101001001","000011001011","101100011110","001010110111","001100000100","101101101001","011111110000","001011101110","000001110011","010111111011","111000100000","011000000010","110100011110","101011011101","100100011111","000110001101","110011100101","011010110101","010001100000","110000110010","111011111001","000000000010","100101010101","110010000110","100001010011","000111110011","111000111111","100011000111","010100111001","001111010010","010111010011","010100001010","111011101101","110000010101","100010010111","101111000111","001100111010","111100110101","011010110010","100010100101","001011011001","010010101111","011101100001","111110101100","100110101001","101110010101","011110101100","001001101000","101100101011","010100100000","011001011001","000110011010","101011000101","010011101000","000000000100","110111000001","011010111110","110001110111","101110111011","101010111001","100111011110","010101101110","010110110000","111001111001","110000000111","010100100001","000100010101","011100101010","100000110100","111000111001","100011100111","111100010111","011001010000","111101111001","101010110110","100100001001","101101111001","110010101010","101110011100","010110111011","100110101011","001101010011","101111001110","000111101010","100000110001","100101110111","000100010000","101110010001","111101011110","111110000001","001001100101","000010011011","010110000010","001001000100","101101011000","110000110110","000000111110","000011000001","010001111010","001100100001","000010010010","010101111111","001010101011","111111000010","111110011000","000010000000","001111000001","101000011110","011010011111","110100100101","100001101000","111100111111","101110110011","100001010001","110001001011","100110111100","010011000000","011010010101","001110000101","001010111001","101010001001","101111011000","110110010111","000100010100","000011000111","110110000100","000000101111","000101001011","101110000001","101011010110","011010011001","100111111001","010111101101","011000011011","000101000010","110000001101","000010010000","000100011000","001001111100","110010000111","001111010110","010110000110","111111100110","001100101111","011111011101","101010101110","000010110111","010011000111","101001101100","001100111000","010110111010","110011111001","100100000110","010110010001","101101001010","101111000001","000100001011","111000111101","100101000001","001110011000","011010101011","101001110010","110110010010","110111110000","011001001101","111001010000","110100011100","110001010101","110010010011","110000111000","000101011011","110100111001","100011110111","101010100101","110100111011","110111001011","010111000100","101000011000","011100010000","111111100000","010100111101","110101010100","011001110101","010000100110","000000001010","000111000101","101000011010","000110010001","110100000011","000001001101","101000100101","101011100011","110110101001","001101001110","000111000110","010011100101","100110010011","001101000011","010010010000","110011010110","101000001100","011011011111","100001100110","010100101100","010110000101","110111111111","101100111000","010110010010","100100100011","010111100111","100000100011","110011001101","000111010001","001001111110","000111010100","000111100100","011110011010","111111100100","110101001010","000110000101","011011111001","100011011101","100110100111","010101001111","110000110000","001000000000","000100011111","111001100101","000110001011","001101010101","110000101001","001100010010","100000111011","100111000000","110000000110","001100001011","100110110011","001001110100","000010011101","000100001010","001111010000","111110100010","011011100111","001101001001","110101000100","011000101111","010001110101","000000011001","010000110101","001001100011","111001000111","000000010010","101110111000","001110001100","000000000101","101011011011","000110010000","000111001100","011101010010","100010011101","100101011001","011010000100","110101110100","001101000101","101101010000","100010111110","001000011001","011110100001","000110010111","101110100111","110001000001","111101100110","110001101000","011001101100","110011011000","011010011100","011110010101","111010101001","111110000101","010111100000","111110001000","011101111100","011011000110","111100011000","001000000001","010011101010","001011111011","011000100001","001101000100","101011001101","110010010000","100000001111","110110100000","001010101101","010000111010","011101100111","000101111000","001110001000","011010111010","101110011011","101000100001","001010001001","101000110101","011111100001","000111110111","110111111011","011011010101","010000111001","101001000001","011001011000","000010000010","111100100011","011111100101","011111001100","100110000000","111110100011","011000000011","101101010001","001011110010","001111010001","000111001011","111110011010","100100111110","011011111000","000111111001","000010010001","000100111010","101011100111","000011001001","100011111111","011100010110","001111011110","010001111101","010100110001","011101000100","101110000000","000011011100","000010010101","011111001000","110000010111","101100010000","111010101110","001010111000","111110011101","100110011111","010001010010","010110110110","000011011010","010000001111","111101100001","001111000110","101100011001","001000100011","010111001001","011111110011","000010110011","000110100111","001000001011","111011110011","011001101110","111101001011","111111110010","000010011111","010000100101","100010111111","101011101111","110001100100","001100110110","100110111101","110110100001","001011101111","000010100011","011101100010","011000110000","010101110010","101010111010","100001000001","100010001011","001110000010","100011101000","101101100000","100111100111","010101010011","101010001111","010111001111","101101000111","000000110101","110000100101","100101000100","000011101101","110011101100","000010010111","100010001111","111010110110","000010100100","110110101000","110011101010","101101001001","110111101000","001101000000","001011100011","110001110001","101000110010","000101110000","011010111111","111000001011","010110101000","011000100100","011100011001","011001010100","010100011010","110110001110","011110000111","101010001010","001000000100","010111110000","101001111111","000101110010","111111001010","011110100100","111110111000","001101001010","000001110000","001111110000","100101010110","111111110011","011011011101","001110010101","111101101110","110100000110","100010000001","101011111101","000110011111","101101010011","100000001110","100100100100","010010111100","000000000000","011111110010","100011100001","100110101111","111011011000","101011001000","111100000110","010000000011","010110011000","010000011001","011011001111","110010101111","111100010101","001111100100","100000011111","000111110000","000101000100","111010100001","000100001111","111100110110","111011101111","101010100010","101100111001","010000001101","111101011000","001011010111","001000101111","111110101101","101100110111","111000010110","110110111101");
	constant expected_output	: word_array := ("010011100111","000110111111","000001110101","110001110101","010011100111","000110110011","111111101111","110111111101","111001010111","110000101101","111010101101","000001110101","010010110111","101010101011","010010010111","101101010101","010010001001","101110111011","110110110001","010111010101","110110000111","101011110111","001001110001","010001011001","101010010111","000111110101","001110100001","101001011101","001101110111","111111100011","001011010111","001001011101","101100111101","010011110001","001000111101","010110111011","001011001111","000011000001","110111111011","011000101011","010100000111","110101111101","111001111001","101011110111","101111101001","110011100111","000110101011","000011000011","010100101011","011000010011","111000010101","000100010001","111111010001","010001101101","000101110111","000110001011","001000110111","111011101101","101100101001","000101101001","000001110101","001110111101","000101001111","000011001011","101101011001","110000000011","110110101101","101101100101","111011010011","010100101001","010001111001","111101000111","010000010011","001001011001","000001101111","111011011111","010110000111","000110010111","111010111101","000000101111","010000000101","101100111111","101011001111","101011101001","010101111101","111001110001","010011101101","001001001101","010000011011","001010011001","000101101011","010011011111","001110000111","101011100111","101000000001","001110100001","000101111101","111000000101","000111011011","000101101101","000110111111","111001010001","010010001011","010010001001","110100100011","010111110111","011000101111","110011111011","000100110011","001110000011","111010011101","010100001111","100111010111","111001110001","000010010101","000111111111","010010110001","111010001001","110010001101","111011110101","101010101111","110100011011","101011000111","010001001111","101111011011","010101101111","110100110111","111000001111","000111000111","101100011011","101011011011","111011100001","101010110101","111100100011","000001100111","101001111001","001000100011","000101111011","100111011101","111011111001","010001101001","101000100111","010110001111","110100100111","110110000001","101110000101","001101100101","111000111111","001110100101","010001000101","110000100011","111101111001","000101010101","101011100011","101000000111","111100100111","010001100111","111001100101","010100000101","110000010101","000111001011","101101100011","110110100111","110100011111","001010001001","010110000101","000101111011","000010011111","100111110001","110111010011","100111111111","111110111111","110000000111","010011101001","111000101111","010100111111","010010010101","001011001001","001111100101","001010011011","110100001011","111001011011","110000001001","010000100011","000000010101","001101001011","000100001011","001000101101","001001100011","110111000001","000001001001","010001101011","001110101011","101111000101","110001001111","110111100101","111110100011","000010011111","000110101111","111011011011","001000110001","111101011011","101100101111","000110000011","010010110111","001000100001","110000010001","101011100001","011001000001","000101111101","101011111011","111010100111","110110000001","111111111101","001110011011","111100100101","110000101011","010100011111","010100111101","111111000101","001010110111","001111100001","001110100011","011000000001","101111010011","010100010111","110110001101","111101101001","101010100011","011001000011","001111111001","101101011111","000110110011","010011111011","111000001001","000110001111","111000000111","101101000011","101001110011","010000010011","000000101101","111100110111","010010101001","101101110101","111001101111","101001110111","111100110111","111100000111","111011011111","100111101011","010011001011","111010011001","111001111101","011001000001","111000001111","001010000101","110111010111","010000011111","100111100001","111010011101","111000111011","001010101101","111011111111","000111100101","011000010111","101111100011","010111110011","010101111101","001010101011","100111100001","101101111111","101100000011","111010111011","011000001001","111010000001","101000101101","111110001101","101101101111","110000101011","110101000111","101100111001","000110111011","101011100011","011000010011","100111001111","010110010111","010111111001","111001100011","010011111011","001101110011","010000011101","011000010011","010101011111","000000111111","110110000001","110111011101","101010011101","010100000111","111000101001","101011101001","111101011011","110111011101","111110101001","000111111011","000100010001","010110000001","101010101011","111001110101","101000101101","000011010101","001101110011","110000001011","001111000111","101100111011","001000010111","101110101101","101011110011","011000011101","101000011001","101000001001","010010110011","010011101011","110101000111","101010010111","111010110011","111010010001","110010100111","001001001011","101010001011","010000011101","110000100001","101110010001","101111111011","001101101001","101101110001","101000100111","110110110111","010111101111","001100010101","001101010101","000101111001","010100010001","000010011101","101001100001","000010110111","001100101001","101011010101","110010100001","101000010011","110011101111","110110110001","101100000011","100110111101","011000110101","010001100101","100111111011","111010000101","111010000101","101110000011","110111111111","001011010101","110000100011","010000110111","101010100011","001001111111","101010011111","111100110001","000111111111","011000011011","101001111111","010010111101","110101000111","000111010001","111110011001","001010100101","010001110101","000000101001","001000100011","101011100111","101000010001","010110100011","000110001111","101101101011","000001010111","001110000001","010011010111","101101101011","001000011111","111001101101","010001100011","101100000111","010010001101","010000110001","101100010001","001010100011","000110001011","110010001001","001011111101","010010111101","000101011101","111001100011","001100111101","101100101101","110000111011","101111010111","001100100100","000101101101","010111001011","001001010011","101010110001","000111100001","111001001101","111011010101","111100101111","010000001001","000000101001","101111101011","010000101001","000101011001","010001110101","110110001001","111100101101","111010000001","110010100011","010010101011","110100000001","110010111011","111000111111","010000110111","100110111111","101101111101","110001001011","110001101111","011000101001","001100011011","110111111101","001000010111","101000110001","110111110001","001000000101","111001010001","111000000011","000100100001","001101001001","110011000001","001000010011","110011110011","111111101111","000000000011","010001111111","010010101011","101010110111","000111000111","010110000101","010100100011","110010100011","111000010011","111001000101","010111101011","010101011101","101101111111","000111010011","010010110111","101110110011","101101101111","110011111111","111111001111","010111111011","101011110011","110100110001","010001101011","010010110111","101110010001","000010010011","010000111001","101110110011","101000100111","101110000101","110010111101","010001100001","000011001101","001111000011","000101111111","111011011011","000110100011","111100110101","000101110001","111111000101","000010010111","000100110101","010100011101","000100000101","100111010111","010011110011","001000111101","000101111111","001011011011","010000101111","010110100101","101011000011","010101001001","010100000011","011001000111","000100000101","110111011011","001011110011","000001111001","001001001001","110000001001","010110100001","000000110001","010011010111","101111000011","111101101001","010110111011","111110000111","010011110011","101101101101","010101001001","010110110011","111010100101","101000000101","101011110001","001111100001","010100011011","111010110101","100111110011","101110101101","110001010011","000101011001","101000110011","010110111101","001011011001","000100010011","110111011101","010101111101","001100000001","111000101111","001101011111","001100110001","011000100011","001110010001","111101011011","010010110111","111100110011","101101010111","110111001011","010110010011","101010100111","000101110111","010100111111","111100000111","111101001101","000000000011","101101111101","101111110011","110010110001","010110000011","101100001101","110100011111","010010111011","001111110111","001010010001","000100101011","101000010011","111000011001","101101001001","111010111111","010101111101","111101101101","000111010011","111001111101","010101100101","000111001011","000111001001","111111101001","110111000111","101101000111","000110011111","001010000101","111010101101","001111011111","000111100011","010101000101","101011111001","000111000001","000000000011","111000011001","000111000101","111100010001","111001100101","110100001001","110111001011","010100010011","010010100101","111101100001","101011110011","001011100111","010111111001","010000111111","110111010011","101001000111","101110011111","101001011011","000111001111","111111011101","110010010011","110010101101","110101110101","101010110101","111001111011","010010111011","101111011111","010010110101","101111000111","010110010011","110000100011","110010010101","000001011001","110100101101","111110110101","111111011111","010010000011","000000110001","010000000101","000011000011","101011011111","101011000001","011000110101","011000000011","001000101001","010100011111","000001011011","000101001101","010110000001","111111101011","101000000101","000000110011","010100100001","110110000001","000110100001","111100110001","110101001101","100111101101","110100010111","110010101011","101100010111","101101000011","010000100101","001001111101","000011101011","000011010101","110010000101","111010000101","111000010011","010111100101","010100010011","110010100001","011000110111","000010010001","111010011111","110011011101","010010010001","110011110101","001111110101","010001111001","010110001011","101010101101","000010110111","000001001001","010110010011","101100110011","010100101001","001111010101","100111001111","000101011001","000111001111","111010101101","000111010111","001100000001","101101011101","010001111101","001001001011","111011101111","110000101001","010011010111","101101000101","110000101011","001011001101","111101111011","110101110111","010100100001","001101000001","111001111001","101100011011","111101101111","001000000001","111110001101","101100001001","101110101111","111010011111","101011100001","000010000001","101010100011","101101010001","101011110101","110100100101","101001110011","001001101101","111001011011","001110010101","111111110111","010011010111","111101010111","001100001011","010011100011","000000000101","000111000001","111000100011","010101011001","110110011011","011000011011","111010110101","110001001111","111100100011","000101001011","000011001001","010100011101","111000111011","001101100101","010001010001","110000010001","110100011011","010000110001","111000100011","001011010001","010000101001","101100111101","111011011101","010000001111","101111001001","010011011011","110101001101","111000101101","010010011011","000110010001","000010100101","001010111101","000111101001","111111101111","101011111001","000011010101","001100100111","110101010001","101111111001","000111001001","110010101101","010110110001","000001111011","111101101011","010100100011","010100101001","111000101101","001100011111","101110011011","110000011001","110001101101","010011110111","101111101101","010100100111","010100010111","011000000001","000101100111","100111011101","010010010101","000100110111","110011110001","000110000011","010011100011","011000100101","010011000111","000010111011","111110010001","000000001001","101111000011","000011111011","000000000001","110000101111","000011000101","010110101011","000110110101","110101100111","101101011111","010001000001","101111110011","010101111111","101101111111","111001001111","010110011001","000110011111","010110101011","110001100011","101100011111","100111101111","111010000011","010000001111","111010001001","001100001001","001010000111","110001100011","111011110101","001001111111","111111010001","001111010101","000111100101","100111111001","010101001111","010010010101","010010010011","001110010011","010101100011","111010110001","101111100001","110110110101","101011001001","000110000001","010010101101","000110001101","000001100111","000111011001","010010101111","101110001001","110110100101","010000101101","101100010111","010001001101","001000110011","111100011111","000110010101","010100010011","111010001001","001001010011","000000100011","100111110111","001110001101","000110110111","110001101101","111110011001","001000011011","111010010011","000101000011","000100110011","000101110001","111111001011","111010010011","001010110111","010110011111","010101001111","000001100111","111011000001","010111000001","110000010111","001101000011","010011110101","000100001001","010001110001","001101001011","111010000111","000001100111","000000110011","010001001111","101010111011","111011010111","101101110001","000011000001","111111100111","110101001011","010001101111","001110011011","000010111001","001010000101","111110101011","000101110101","111011011011","010100111101","001100001001","010000110101","000010001101","010101110101","010110101101","111110100101","000111100001","101010111011","100110111101","010101100111","010100111001","101110100001","111010110001","101011011111","010101001001","110110001101","111101011111","000011100111","000100110011","010010010101","001111100111","010011011101","101100100011","110010110111","111000001101","000011010101","101101000101","110001000111","111010000101","000101011101","101111110011","010100000011","101101011001","000000001111","111100010101","101100101011","000011110001","101011110111","010111100011","110101010001","111011011011","000000101001","111101011101","101111111011","101100110001","110010011101","001011000101","000101001101","111011011001","101100001011","001000100101","001001111001","110101100001","010010100101","010001011011","001100110111","010000001101","000101001011","110100011001","000111001111","110111011011","010010111001","000101010101","110011010001","010000001111","101000001011","010010111111","100111010011","010100010101","010111101111","010101010111","111001110111","111111111011","001100011101","010000111001","111000010011","111011110011","101111000111","111011001001","000010001001","111000001101","110111111101","111001110001","010010100101","000000000000","000111110001","110001001111","110010010101","111110100011","101101000111","100111111101","010101011001","001111110111","010101001101","001101000111","101101101101","111110111001","010011010011","101111110111","000011111001","010000001001","101001011101","000011010011","111110001101","101000110001","111001010001","110111000111","010001111111","101111111011","000111000101","000010110001","111110111001","111010110111","111101011111","101011000011");

begin

	cordicAtan2UnderTest : CORDICAtan2
		port map (
			clock		=> test_clock,
			reset		=> test_reset,
			inA			=> test_inA,
			inB			=> test_inB,
			valid		=> test_valid,
			atan2Out	=> test_output
		);

	test_clock <= (not test_end) and (not test_clock) after 50ns;

	-- stimuli
	driveProcess : process
	begin
		wait for 60ns;
		
		test_reset <= '0';

		for i in 0 to TEST_SIZE-1 loop
			test_inA <= test_inputA(i);
			test_inB <= test_inputB(i);

			for j in 0 to LUT_SIZE-1 loop
				wait until rising_edge(test_clock);
			end loop;

			test_expected <= expected_output(i);

			wait for 25ns;

			if test_valid = '1' and test_output = expected_output(i) then
				test_correct <= '1';
			else
				test_correct <= '0';
			end if;

			assert (test_valid = '1' and test_output = expected_output(i))
			report "ERROR: detected for index i = " & integer'image(i)
				& "; A = " & integer'image(to_integer(signed(test_inA)))
				& "; B = " & integer'image(to_integer(signed(test_inB)))
				& "."
			severity error;

		end loop;

		wait for 100ns;

		test_end <= '1';

		wait;
	end	process;
	
end System_TB_Arch;